module projeto();
endmodule
